module top_module( input in, output out );
	assign out = ~in;     // ~ is bitwise-NOT  and ! is logic-NOT
endmodule
